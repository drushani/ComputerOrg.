/*
	Input Port
		1. immed_in: Ū�J����sign extend���
	Output Port
		1. ext_immed_out: ��X�w����sign extend���
*/
module sign_extend( immed_in, ext_immed );
	input[15:0] immed_in;
	output[31:0] ext_immed;
	assign ext_immed = { {16{immed_in[15]}}, immed_in };
endmodule
