module shifter( dataA, dataB, dataOut );

input [31:0] dataA ;
input [4:0] dataB ;
output [31:0] dataOut ;
wire [31:0] temp0, temp1, temp2, temp3, temp4 ;

// 1
mux2_1 m1_1(dataB[0], dataA[1], dataA[0], temp0[0]);
mux2_1 m1_2(dataB[0], dataA[2], dataA[1], temp0[1]);
mux2_1 m1_3(dataB[0], dataA[3], dataA[2], temp0[2]);
mux2_1 m1_4(dataB[0], dataA[4], dataA[3], temp0[3]);
mux2_1 m1_5(dataB[0], dataA[5], dataA[4], temp0[4]);
mux2_1 m1_6(dataB[0], dataA[6], dataA[5], temp0[5]);
mux2_1 m1_7(dataB[0], dataA[7], dataA[6], temp0[6]);
mux2_1 m1_8(dataB[0], dataA[8], dataA[7], temp0[7]);
mux2_1 m1_9(dataB[0], dataA[9], dataA[8], temp0[8]);
mux2_1 m1_10(dataB[0], dataA[10], dataA[9], temp0[9]);
mux2_1 m1_11(dataB[0], dataA[11], dataA[10], temp0[10]);
mux2_1 m1_12(dataB[0], dataA[12], dataA[11], temp0[11]);
mux2_1 m1_13(dataB[0], dataA[13], dataA[12], temp0[12]);
mux2_1 m1_14(dataB[0], dataA[14], dataA[13], temp0[13]);
mux2_1 m1_15(dataB[0], dataA[15], dataA[14], temp0[14]);
mux2_1 m1_16(dataB[0], dataA[16], dataA[15], temp0[15]);
mux2_1 m1_17(dataB[0], dataA[17], dataA[16], temp0[16]);
mux2_1 m1_18(dataB[0], dataA[18], dataA[17], temp0[17]);
mux2_1 m1_19(dataB[0], dataA[19], dataA[18], temp0[18]);
mux2_1 m1_20(dataB[0], dataA[20], dataA[19], temp0[19]);
mux2_1 m1_21(dataB[0], dataA[21], dataA[20], temp0[20]);
mux2_1 m1_22(dataB[0], dataA[22], dataA[21], temp0[21]);
mux2_1 m1_23(dataB[0], dataA[23], dataA[22], temp0[22]);
mux2_1 m1_24(dataB[0], dataA[24], dataA[23], temp0[23]);
mux2_1 m1_25(dataB[0], dataA[25], dataA[24], temp0[24]);
mux2_1 m1_26(dataB[0], dataA[26], dataA[25], temp0[25]);
mux2_1 m1_27(dataB[0], dataA[27], dataA[26], temp0[26]);
mux2_1 m1_28(dataB[0], dataA[28], dataA[27], temp0[27]);
mux2_1 m1_29(dataB[0], dataA[29], dataA[28], temp0[28]);
mux2_1 m1_30(dataB[0], dataA[30], dataA[29], temp0[29]);
mux2_1 m1_31(dataB[0], dataA[31], dataA[30], temp0[30]);
mux2_1 m1_32(dataB[0], 1'b0, dataA[31], temp0[31]);

// 2
mux2_1 m2_1(dataB[1], temp0[2], temp0[0], temp1[0]);
mux2_1 m2_2(dataB[1], temp0[3], temp0[1], temp1[1]);
mux2_1 m2_3(dataB[1], temp0[4], temp0[2], temp1[2]);
mux2_1 m2_4(dataB[1], temp0[5], temp0[3], temp1[3]);
mux2_1 m2_5(dataB[1], temp0[6], temp0[4], temp1[4]);
mux2_1 m2_6(dataB[1], temp0[7], temp0[5], temp1[5]);
mux2_1 m2_7(dataB[1], temp0[8], temp0[6], temp1[6]);
mux2_1 m2_8(dataB[1], temp0[9], temp0[7], temp1[7]);
mux2_1 m2_9(dataB[1], temp0[10], temp0[8], temp1[8]);
mux2_1 m2_10(dataB[1], temp0[11], temp0[9], temp1[9]);
mux2_1 m2_11(dataB[1], temp0[12], temp0[10], temp1[10]);
mux2_1 m2_12(dataB[1], temp0[13], temp0[11], temp1[11]);
mux2_1 m2_13(dataB[1], temp0[14], temp0[12], temp1[12]);
mux2_1 m2_14(dataB[1], temp0[15], temp0[13], temp1[13]);
mux2_1 m2_15(dataB[1], temp0[16], temp0[14], temp1[14]);
mux2_1 m2_16(dataB[1], temp0[17], temp0[15], temp1[15]);
mux2_1 m2_17(dataB[1], temp0[18], temp0[16], temp1[16]);
mux2_1 m2_18(dataB[1], temp0[19], temp0[17], temp1[17]);
mux2_1 m2_19(dataB[1], temp0[20], temp0[18], temp1[18]);
mux2_1 m2_20(dataB[1], temp0[21], temp0[19], temp1[19]);
mux2_1 m2_21(dataB[1], temp0[22], temp0[20], temp1[20]);
mux2_1 m2_22(dataB[1], temp0[23], temp0[21], temp1[21]);
mux2_1 m2_23(dataB[1], temp0[24], temp0[22], temp1[22]);
mux2_1 m2_24(dataB[1], temp0[25], temp0[23], temp1[23]) ;
mux2_1 m2_25(dataB[1], temp0[26], temp0[24], temp1[24]) ;
mux2_1 m2_26(dataB[1], temp0[27], temp0[25], temp1[25]) ;
mux2_1 m2_27(dataB[1], temp0[28], temp0[26], temp1[26]) ;
mux2_1 m2_28(dataB[1], temp0[29], temp0[27], temp1[27]) ;
mux2_1 m2_29(dataB[1], temp0[30], temp0[28], temp1[28]) ;
mux2_1 m2_30(dataB[1], temp0[31], temp0[29], temp1[29]) ;
mux2_1 m2_31(dataB[1], 1'b0, temp0[30], temp1[30]) ;
mux2_1 m2_32(dataB[1], 1'b0, temp0[31], temp1[31]) ;

// 4
mux2_1 m3_1(dataB[2], temp1[4], temp1[0], temp2[0]);
mux2_1 m3_2(dataB[2], temp1[5], temp1[1], temp2[1]);
mux2_1 m3_3(dataB[2], temp1[6], temp1[2], temp2[2]);
mux2_1 m3_4(dataB[2], temp1[7], temp1[3], temp2[3]);
mux2_1 m3_5(dataB[2], temp1[8], temp1[4], temp2[4]);
mux2_1 m3_6(dataB[2], temp1[9], temp1[5], temp2[5]);
mux2_1 m3_7(dataB[2], temp1[10], temp1[6], temp2[6]);
mux2_1 m3_8(dataB[2], temp1[11], temp1[7], temp2[7]);
mux2_1 m3_9(dataB[2], temp1[12], temp1[8], temp2[8]);
mux2_1 m3_10(dataB[2], temp1[13], temp1[9], temp2[9]);
mux2_1 m3_11(dataB[2], temp1[14], temp1[10], temp2[10]);
mux2_1 m3_12(dataB[2], temp1[15], temp1[11], temp2[11]);
mux2_1 m3_13(dataB[2], temp1[16], temp1[12], temp2[12]);
mux2_1 m3_14(dataB[2], temp1[17], temp1[13], temp2[13]);
mux2_1 m3_15(dataB[2], temp1[18], temp1[14], temp2[14]);
mux2_1 m3_16(dataB[2], temp1[19], temp1[15], temp2[15]);
mux2_1 m3_17(dataB[2], temp1[20], temp1[16], temp2[16]);
mux2_1 m3_18(dataB[2], temp1[21], temp1[17], temp2[17]);
mux2_1 m3_19(dataB[2], temp1[22], temp1[18], temp2[18]);
mux2_1 m3_20(dataB[2], temp1[23], temp1[19], temp2[19]);
mux2_1 m3_21(dataB[2], temp1[24], temp1[20], temp2[20]);
mux2_1 m3_22(dataB[2], temp1[25], temp1[21], temp2[21]);
mux2_1 m3_23(dataB[2], temp1[26], temp1[22], temp2[22]);
mux2_1 m3_24(dataB[2], temp1[27], temp1[23], temp2[23]);
mux2_1 m3_25(dataB[2], temp1[28], temp1[24], temp2[24]);
mux2_1 m3_26(dataB[2], temp1[29], temp1[25], temp2[25]);
mux2_1 m3_27(dataB[2], temp1[30], temp1[26], temp2[26]);
mux2_1 m3_28(dataB[2], temp1[31], temp1[27], temp2[27]);
mux2_1 m3_29(dataB[2], 1'b0, temp1[28], temp2[28]);
mux2_1 m3_30(dataB[2], 1'b0, temp1[29], temp2[29]);
mux2_1 m3_31(dataB[2], 1'b0, temp1[30], temp2[30]);
mux2_1 m3_32(dataB[2], 1'b0, temp1[31], temp2[31]);

// 8
mux2_1 m4_1(dataB[3], temp2[8], temp2[0], temp3[0]);
mux2_1 m4_2(dataB[3], temp2[9], temp2[1], temp3[1]);
mux2_1 m4_3(dataB[3], temp2[10], temp2[2], temp3[2]);
mux2_1 m4_4(dataB[3], temp2[11], temp2[3], temp3[3]);
mux2_1 m4_5(dataB[3], temp2[12], temp2[4], temp3[4]);
mux2_1 m4_6(dataB[3], temp2[13], temp2[5], temp3[5]);
mux2_1 m4_7(dataB[3], temp2[14], temp2[6], temp3[6]);
mux2_1 m4_8(dataB[3], temp2[15], temp2[7], temp3[7]);
mux2_1 m4_9(dataB[3], temp2[16], temp2[8], temp3[8]);
mux2_1 m4_10(dataB[3], temp2[17], temp2[9], temp3[9]);
mux2_1 m4_11(dataB[3], temp2[18], temp2[10], temp3[10]);
mux2_1 m4_12(dataB[3], temp2[19], temp2[11], temp3[11]);
mux2_1 m4_13(dataB[3], temp2[20], temp2[12], temp3[12]);
mux2_1 m4_14(dataB[3], temp2[21], temp2[13], temp3[13]);
mux2_1 m4_15(dataB[3], temp2[22], temp2[14], temp3[14]);
mux2_1 m4_16(dataB[3], temp2[23], temp2[15], temp3[15]);
mux2_1 m4_17(dataB[3], temp2[24], temp2[16], temp3[16]);
mux2_1 m4_18(dataB[3], temp2[25], temp2[17], temp3[17]);
mux2_1 m4_19(dataB[3], temp2[26], temp2[18], temp3[18]);
mux2_1 m4_20(dataB[3], temp2[27], temp2[19], temp3[19]);
mux2_1 m4_21(dataB[3], temp2[28], temp2[20], temp3[20]);
mux2_1 m4_22(dataB[3], temp2[29], temp2[21], temp3[21]);
mux2_1 m4_23(dataB[3], temp2[30], temp2[22], temp3[22]);
mux2_1 m4_24(dataB[3], temp2[31], temp2[23], temp3[23]);
mux2_1 m4_25(dataB[3], 1'b0, temp2[24], temp3[24] ) ;
mux2_1 m4_26(dataB[3], 1'b0, temp2[25], temp3[25] ) ;
mux2_1 m4_27(dataB[3], 1'b0, temp2[26], temp3[26] ) ;
mux2_1 m4_28(dataB[3], 1'b0, temp2[27], temp3[27] ) ;
mux2_1 m4_29(dataB[3], 1'b0, temp2[28], temp3[28] ) ;
mux2_1 m4_30(dataB[3], 1'b0, temp2[29], temp3[29] ) ;
mux2_1 m4_31(dataB[3], 1'b0, temp2[30], temp3[30] ) ;
mux2_1 m4_32(dataB[3], 1'b0, temp2[31], temp3[31] ) ;

// 16
mux2_1 m5_1(dataB[4], temp3[16], temp3[0], temp4[0]);
mux2_1 m5_2(dataB[4], temp3[17], temp3[1], temp4[1]);
mux2_1 m5_3(dataB[4], temp3[18], temp3[2], temp4[2]);
mux2_1 m5_4(dataB[4], temp3[19], temp3[3], temp4[3]);
mux2_1 m5_5(dataB[4], temp3[20], temp3[4], temp4[4]);
mux2_1 m5_6(dataB[4], temp3[21], temp3[5], temp4[5]);
mux2_1 m5_7(dataB[4], temp3[22], temp3[6], temp4[6]);
mux2_1 m5_8(dataB[4], temp3[23], temp3[7], temp4[7]);
mux2_1 m5_9(dataB[4], temp3[24], temp3[8], temp4[8]);
mux2_1 m5_10(dataB[4], temp3[25], temp3[9], temp4[9]);
mux2_1 m5_11(dataB[4], temp3[26], temp3[10], temp4[10]);
mux2_1 m5_12(dataB[4], temp3[27], temp3[11], temp4[11]);
mux2_1 m5_13(dataB[4], temp3[28], temp3[12], temp4[12]);
mux2_1 m5_14(dataB[4], temp3[29], temp3[13], temp4[13]);
mux2_1 m5_15(dataB[4], temp3[30], temp3[14], temp4[14]);
mux2_1 m5_16(dataB[4], temp3[31], temp3[15], temp4[15]);
mux2_1 m5_17(dataB[4], 1'b0, temp3[16], temp4[16]);
mux2_1 m5_18(dataB[4], 1'b0, temp3[17], temp4[17]);
mux2_1 m5_19(dataB[4], 1'b0, temp3[18], temp4[18]);
mux2_1 m5_20(dataB[4], 1'b0, temp3[19], temp4[19]);
mux2_1 m5_21(dataB[4], 1'b0, temp3[20], temp4[20]);
mux2_1 m5_22(dataB[4], 1'b0, temp3[21], temp4[21]);
mux2_1 m5_23(dataB[4], 1'b0, temp3[22], temp4[22]);
mux2_1 m5_24(dataB[4], 1'b0, temp3[23], temp4[23]);
mux2_1 m5_25(dataB[4], 1'b0, temp3[24], temp4[24]);
mux2_1 m5_26(dataB[4], 1'b0, temp3[25], temp4[25]);
mux2_1 m5_27(dataB[4], 1'b0, temp3[26], temp4[26]);
mux2_1 m5_28(dataB[4], 1'b0, temp3[27], temp4[27]);
mux2_1 m5_29(dataB[4], 1'b0, temp3[28], temp4[28]);
mux2_1 m5_30(dataB[4], 1'b0, temp3[29], temp4[29]);
mux2_1 m5_31(dataB[4], 1'b0, temp3[30], temp4[30]);
mux2_1 m5_32(dataB[4], 1'b0, temp3[31], temp4[31]);

assign dataOut = temp4 ; 

endmodule